        bins pos0             = {128'h00000000000000000000000000000000};
        bins neg0             = {128'h80000000000000000000000000000000};
        bins pos1             = {128'h3FFF0000000000000000000000000000};
        bins neg1             = {128'hBFFF0000000000000000000000000000};
        bins pos1p5           = {128'h3FFF8000000000000000000000000000};
        bins neg1p5           = {128'hBFFF8000000000000000000000000000};
        bins pos2             = {128'h40000000000000000000000000000000};
        bins neg2             = {128'hc0000000000000000000000000000000};
        bins posminnorm       = {128'h00010000000000000000000000000000};
        bins negminnorm       = {128'h80010000000000000000000000000000};
        bins posmaxnorm       = {128'h7FFEFFFFFFFFFFFFFFFFFFFFFFFFFFFF};
        bins negmaxnorm       = {128'hFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFF};
        // bins posnorm          = {[128'h00010000000000000000000000000001:128'h7FFEFFFFFFFFFFFFFFFFFFFFFFFFFFFE]};
        // bins negnorm          = {[128'h80010000000000000000000000000001:128'hFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFE]};
        bins posmax_subnorm   = {128'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFF};
        bins negmax_subnorm   = {128'h8000FFFFFFFFFFFFFFFFFFFFFFFFFFFF};
        // bins posmid_subnorm   = {128'h0000E000000000000000000000000000};
        // bins negmid_subnorm   = {128'h8000E000000000000000000000000000};
        bins posmin_subnorm   = {128'h00000000000000000000000000000001};
        bins negmin_subnorm   = {128'h80000000000000000000000000000001};
        bins pos_subnorm      = {[128'h00000000000000000000000000000002:128'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFE]};
        bins neg_subnorm      = {[128'h80000000000000000000000000000002:128'h8000FFFFFFFFFFFFFFFFFFFFFFFFFFFE]};  
        bins posinfinity      = {128'h7FFF0000000000000000000000000000};
        bins neginfinity      = {128'hFFFF0000000000000000000000000000};
        bins posQNaN          = {[128'h7FFF8000000000000000000000000000:128'h7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF]};
        bins posSNaN          = {[128'h7FFF0000000000000000000000000001:128'h7FFF7FFFFFFFFFFFFFFFFFFFFFFFFFFF]};
        bins negQNaN          = {[128'hFFFF8000000000000000000000000000:128'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF]};
        bins negSNaN          = {[128'hFFFF0000000000000000000000000001:128'hFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFF]};
