        // all conversion operations
        bins op_cfi    = {[OP_CFI  : OP_CFI  | 32'hF]};
        bins op_cff    = {[OP_CFF   : OP_CFF   | 32'hF]}; 