        bins pos0             = {16'h0000};
        bins neg0             = {16'h8000};
        bins pos1             = {16'h3f80};
        bins neg1             = {16'hbf80};
        bins pos1p5           = {16'h3fc0};
        bins neg1p5           = {16'hbfc0};
        bins pos2             = {16'h4000};
        bins neg2             = {16'hc000};
        bins posminnorm       = {16'h0080};
        bins negminnorm       = {16'h8080};
        bins posmaxnorm       = {16'h7f7f};
        bins negmaxnorm       = {16'hff7f};
        bins posnorm          = {[16'h0081:16'h7f7e]};
        bins negnorm          = {[16'h8081:16'hff7e]};
        bins posmax_subnorm   = {16'h007f};
        bins negmax_subnorm   = {16'h807f};
        // bins posmid_subnorm   = {16'h0040};
        // bins negmid_subnorm   = {16'h8040};
        bins posmin_subnorm   = {16'h0001};
        bins negmin_subnorm   = {16'h8001};
        bins pos_subnorm      = {[16'h0002:16'h007e]};
        bins neg_subnorm      = {[16'h8002:16'h807e]};
        bins posinfinity      = {16'h7f80};
        bins neginfinity      = {16'hff80};
        `ifndef IGNORE_NANS
            bins posQNaN          = {[16'h7fc0:16'h7fff]};
            bins posSNaN          = {[16'h7f81:16'h7fbf]};
            bins negQNaN          = {[16'hffc0:16'hffff]};
            bins negSNaN          = {[16'hff81:16'hffbf]};
        `endif
