// define macros for which models to check coverage for
// e.g. `define COVER_B1 for model B1

`define COVER_B1
// `define COVER_B2
// `define COVER_B3
// `define COVER_B4
// `define COVER_B5
// `define COVER_B6
// `define COVER_B7
// `define COVER_B8
`define COVER_B9
`define COVER_B10
// `define COVER_B11
`define COVER_B12
// `define COVER_B13
`define COVER_B14
// `define COVER_B15
// `define COVER_B16
// `define COVER_B17
// `define COVER_B18
// `define COVER_B19
// `define COVER_B20
`define COVER_B21
// `define COVER_B22
// `define COVER_B23
// `define COVER_B24
// `define COVER_B25
// `define COVER_B26
// `define COVER_B27
// `define COVER_B28
// `define COVER_B29

// define macros for which precisions to check coverage for
// e.g. `define COVER_F32 for single precision

`define COVER_F32
`define COVER_F64
`define COVER_F128
`define COVER_F16
`define COVER_BF16

// define macro for long int support (i.e. 64 bit DUT)

`define COVER_LONG